/* http://srecord.sourceforge.net/ */
@00000000 00200E13 00000093 00000113 0020F663 35C01263 01C01663 FE20FEE3
@00000007 33C01C63 00300E13 00100093 00100113 0020F663 33C01263 01C01663
@0000000E FE20FEE3 31C01C63 00400E13 FFF00093 FFF00113 0020F663 31C01263
@00000015 01C01663 FE20FEE3 2FC01C63 00500E13 00100093 00000113 0020F663
@0000001C 2FC01263 01C01663 FE20FEE3 2DC01C63 00600E13 FFF00093 FFE00113
@00000023 0020F663 2DC01263 01C01663 FE20FEE3 2BC01C63 00700E13 FFF00093
@0000002A 00000113 0020F663 2BC01263 01C01663 FE20FEE3 29C01C63 00800E13
@00000031 00000093 00100113 0020F463 01C01463 29C01063 FE20FEE3 00900E13
@00000038 FFE00093 FFF00113 0020F463 01C01463 27C01263 FE20FEE3 00A00E13
@0000003F 00000093 FFF00113 0020F463 01C01463 25C01463 FE20FEE3 00B00E13
@00000046 800000B7 FFF08093 80000137 0020F463 01C01463 23C01463 FE20FEE3
@0000004D 00C00E13 00000213 F00000B7 FFF08093 F0000137 2020F663 00120213
@00000054 00200293 FE5214E3 00D00E13 00000213 F00000B7 FFF08093 F0000137
@0000005B 00000013 1E20F263 00120213 00200293 FE5212E3 00E00E13 00000213
@00000062 F00000B7 FFF08093 F0000137 00000013 00000013 1A20FC63 00120213
@00000069 00200293 FE5210E3 00F00E13 00000213 F00000B7 FFF08093 00000013
@00000070 F0000137 1820F863 00120213 00200293 FE5212E3 01000E13 00000213
@00000077 F00000B7 FFF08093 00000013 F0000137 00000013 1620F263 00120213
@0000007E 00200293 FE5210E3 01100E13 00000213 F00000B7 FFF08093 00000013
@00000085 00000013 F0000137 1220FC63 00120213 00200293 FE5210E3 01200E13
@0000008C 00000213 F00000B7 FFF08093 F0000137 1020FA63 00120213 00200293
@00000093 FE5214E3 01300E13 00000213 F00000B7 FFF08093 F0000137 00000013
@0000009A 0E20F663 00120213 00200293 FE5212E3 01400E13 00000213 F00000B7
@000000A1 FFF08093 F0000137 00000013 00000013 0C20F063 00120213 00200293
@000000A8 FE5210E3 01500E13 00000213 F00000B7 FFF08093 00000013 F0000137
@000000AF 0820FC63 00120213 00200293 FE5212E3 01600E13 00000213 F00000B7
@000000B6 FFF08093 00000013 F0000137 00000013 0620F663 00120213 00200293
@000000BD FE5210E3 01700E13 00000213 F00000B7 FFF08093 00000013 00000013
@000000C4 F0000137 0420F063 00120213 00200293 FE5210E3 00100093 0000FA63
@000000CB 00108093 00108093 00108093 00108093 00108093 00108093 00300E93
@000000D2 01800E13 01D09463 01C01A63 FF000513 00000593 00B52023 FF5FF06F
@000000D9 FF000513 00100593 00B52023 FF5FF06F
