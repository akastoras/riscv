/* http://srecord.sourceforge.net/ */
@00000000 00200E13 00000093 00100113 0020C663 2BC01863 01C01663 FE20CEE3
@00000007 2BC01263 00300E13 FFF00093 00100113 0020C663 29C01863 01C01663
@0000000E FE20CEE3 29C01263 00400E13 FFE00093 FFF00113 0020C663 27C01863
@00000015 01C01663 FE20CEE3 27C01263 00500E13 00100093 00000113 0020C463
@0000001C 01C01463 25C01663 FE20CEE3 00600E13 00100093 FFF00113 0020C463
@00000023 01C01463 23C01863 FE20CEE3 00700E13 FFF00093 FFE00113 0020C463
@0000002A 01C01463 21C01A63 FE20CEE3 00800E13 00100093 FFE00113 0020C463
@00000031 01C01463 1FC01C63 FE20CEE3 00900E13 00000213 00000093 FFF00113
@00000038 1E20C063 00120213 00200293 FE5216E3 00A00E13 00000213 00000093
@0000003F FFF00113 00000013 1A20CE63 00120213 00200293 FE5214E3 00B00E13
@00000046 00000213 00000093 FFF00113 00000013 00000013 1820CA63 00120213
@0000004D 00200293 FE5212E3 00C00E13 00000213 00000093 00000013 FFF00113
@00000054 1620C863 00120213 00200293 FE5214E3 00D00E13 00000213 00000093
@0000005B 00000013 FFF00113 00000013 1420C463 00120213 00200293 FE5212E3
@00000062 00E00E13 00000213 00000093 00000013 00000013 FFF00113 1220C063
@00000069 00120213 00200293 FE5212E3 00F00E13 00000213 00000093 FFF00113
@00000070 1020C063 00120213 00200293 FE5216E3 01000E13 00000213 00000093
@00000077 FFF00113 00000013 0C20CE63 00120213 00200293 FE5214E3 01100E13
@0000007E 00000213 00000093 FFF00113 00000013 00000013 0A20CA63 00120213
@00000085 00200293 FE5212E3 01200E13 00000213 00000093 00000013 FFF00113
@0000008C 0820C863 00120213 00200293 FE5214E3 01300E13 00000213 00000093
@00000093 00000013 FFF00113 00000013 0620C463 00120213 00200293 FE5212E3
@0000009A 01400E13 00000213 00000093 00000013 00000013 FFF00113 0420C063
@000000A1 00120213 00200293 FE5212E3 00100093 00104A63 00108093 00108093
@000000A8 00108093 00108093 00108093 00108093 00300E93 01500E13 01D09463
@000000AF 01C01A63 FF000513 00000593 00B52023 FF5FF06F FF000513 00100593
@000000B6 00B52023 FF5FF06F
