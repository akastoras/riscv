/* http://srecord.sourceforge.net/ */
@00000000 00200E13 00000093 0100026F 00000013 00000013 0400006F 00000117
@00000007 FF410113 02411A63 00100093 0140006F 00108093 00108093 00108093
@0000000E 00108093 00108093 00108093 00300E93 00300E13 01D09463 01C01A63
@00000015 FF000513 00000593 00B52023 FF5FF06F FF000513 00100593 00B52023
@0000001C FF5FF06F
