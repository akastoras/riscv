/* http://srecord.sourceforge.net/ */
@00000000 000000B7 00000E93 00200E13 05D09A63 FFFFF0B7 4010D093 80000E93
@00000007 00300E13 05D09063 7FFFF0B7 4140D093 7FF00E93 00400E13 03D09663
@0000000E 800000B7 4140D093 80000E93 00500E13 01D09C63 80000037 00000E93
@00000015 00600E13 01D01463 01C01A63 FF000513 00000593 00B52023 FF5FF06F
@0000001C FF000513 00100593 00B52023 FF5FF06F
