/* http://srecord.sourceforge.net/ */
@00000000 00000093 00000113 0020A1B3 00000E93 00200E13 4BD19A63 00100093
@00000007 00100113 0020A1B3 00000E93 00300E13 49D19E63 00300093 00700113
@0000000E 0020A1B3 00100E93 00400E13 49D19263 00700093 00300113 0020A1B3
@00000015 00000E93 00500E13 47D19663 00000093 FFFF8137 0020A1B3 00000E93
@0000001C 00600E13 45D19A63 800000B7 00000113 0020A1B3 00100E93 00700E13
@00000023 43D19E63 800000B7 FFFF8137 0020A1B3 00100E93 00800E13 43D19263
@0000002A 00000093 00008137 FFF10113 0020A1B3 00100E93 00900E13 41D19463
@00000031 800000B7 FFF08093 00000113 0020A1B3 00000E93 00A00E13 3FD19663
@00000038 800000B7 FFF08093 00008137 FFF10113 0020A1B3 00000E93 00B00E13
@0000003F 3DD19663 800000B7 00008137 FFF10113 0020A1B3 00100E93 00C00E13
@00000046 3BD19863 800000B7 FFF08093 FFFF8137 0020A1B3 00000E93 00D00E13
@0000004D 39D19A63 00000093 FFF00113 0020A1B3 00000E93 00E00E13 37D19E63
@00000054 FFF00093 00100113 0020A1B3 00100E93 00F00E13 37D19263 FFF00093
@0000005B FFF00113 0020A1B3 00000E93 01000E13 35D19663 00E00093 00D00113
@00000062 0020A0B3 00000E93 01100E13 33D09A63 00B00093 00D00113 0020A133
@00000069 00100E93 01200E13 31D11E63 00D00093 0010A0B3 00000E93 01300E13
@00000070 31D09463 00000213 00B00093 00D00113 0020A1B3 00018313 00120213
@00000077 00200293 FE5214E3 00100E93 01400E13 2DD31E63 00000213 00E00093
@0000007E 00D00113 0020A1B3 00000013 00018313 00120213 00200293 FE5212E3
@00000085 00000E93 01500E13 2BD31663 00000213 00C00093 00D00113 0020A1B3
@0000008C 00000013 00000013 00018313 00120213 00200293 FE5210E3 00100E93
@00000093 01600E13 27D31C63 00000213 00E00093 00D00113 0020A1B3 00120213
@0000009A 00200293 FE5216E3 00000E93 01700E13 25D19863 00000213 00B00093
@000000A1 00D00113 00000013 0020A1B3 00120213 00200293 FE5214E3 00100E93
@000000A8 01800E13 23D19263 00000213 00F00093 00D00113 00000013 00000013
@000000AF 0020A1B3 00120213 00200293 FE5212E3 00000E93 01900E13 1FD19A63
@000000B6 00000213 00A00093 00000013 00D00113 0020A1B3 00120213 00200293
@000000BD FE5214E3 00100E93 01A00E13 1DD19463 00000213 01000093 00000013
@000000C4 00D00113 00000013 0020A1B3 00120213 00200293 FE5212E3 00000E93
@000000CB 01B00E13 19D19C63 00000213 00900093 00000013 00000013 00D00113
@000000D2 0020A1B3 00120213 00200293 FE5212E3 00100E93 01C00E13 17D19463
@000000D9 00000213 00D00113 01100093 0020A1B3 00120213 00200293 FE5216E3
@000000E0 00000E93 01D00E13 15D19063 00000213 00D00113 00800093 00000013
@000000E7 0020A1B3 00120213 00200293 FE5214E3 00100E93 01E00E13 11D19A63
@000000EE 00000213 00D00113 01200093 00000013 00000013 0020A1B3 00120213
@000000F5 00200293 FE5212E3 00000E93 01F00E13 0FD19263 00000213 00D00113
@000000FC 00000013 00700093 0020A1B3 00120213 00200293 FE5214E3 00100E93
@00000103 02000E13 0BD19C63 00000213 00D00113 00000013 01300093 00000013
@0000010A 0020A1B3 00120213 00200293 FE5212E3 00000E93 02100E13 09D19463
@00000111 00000213 00D00113 00000013 00000013 00600093 0020A1B3 00120213
@00000118 00200293 FE5212E3 00100E93 02200E13 05D19C63 FFF00093 00102133
@0000011F 00000E93 02300E13 05D11263 FFF00093 0000A133 00100E93 02400E13
@00000126 03D11863 000020B3 00000E93 02500E13 03D09063 01000093 01E00113
@0000012D 0020A033 00000E93 02600E13 01D01463 01C01A63 FF000513 00000593
@00000134 00B52023 FF5FF06F FF000513 00100593 00B52023 FF5FF06F
