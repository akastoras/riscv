/* http://srecord.sourceforge.net/ */
@00000000 7FC00097 00008093 00009183 0FF00E93 00200E13 25D19C63 7FC00097
@00000007 FE808093 00209183 F0000E93 00300E13 25D19063 7FC00097 FD008093
@0000000E 00409183 00001EB7 FF0E8E93 00400E13 23D19263 7FC00097 FB408093
@00000015 00609183 FFFFFEB7 00FE8E93 00500E13 21D19463 7FC00097 F9E08093
@0000001C FFA09183 0FF00E93 00600E13 1FD19863 7FC00097 F8608093 FFC09183
@00000023 F0000E93 00700E13 1DD19C63 7FC00097 F6E08093 FFE09183 00001EB7
@0000002A FF0E8E93 00800E13 1BD19E63 7FC00097 F5208093 00009183 FFFFFEB7
@00000031 00FE8E93 00900E13 1BD19063 7FC00097 F3008093 FE008093 02009283
@00000038 0FF00E93 00A00E13 19D29263 7FC00097 F1408093 FFB08093 00709283
@0000003F F0000E93 00B00E13 17D29463 00C00E13 00000213 7FC00097 EF208093
@00000046 00209183 00018313 00001EB7 FF0E8E93 15D31263 00120213 00200293
@0000004D FC521EE3 00D00E13 00000213 7FC00097 EC408093 00209183 00000013
@00000054 00018313 FFFFFEB7 00FE8E93 11D31863 00120213 00200293 FC521CE3
@0000005B 00E00E13 00000213 7FC00097 E8C08093 00209183 00000013 00000013
@00000062 00018313 F0000E93 0DD31E63 00120213 00200293 FC521CE3 00F00E13
@00000069 00000213 7FC00097 E5A08093 00209183 00001EB7 FF0E8E93 0BD19863
@00000070 00120213 00200293 FE5210E3 01000E13 00000213 7FC00097 E3008093
@00000077 00000013 00209183 FFFFFEB7 00FE8E93 09D19063 00120213 00200293
@0000007E FC521EE3 01100E13 00000213 7FC00097 DFC08093 00000013 00000013
@00000085 00209183 F0000E93 05D19863 00120213 00200293 FC521EE3 7FC00297
@0000008C DD428293 00029103 00200113 00200E93 01200E13 03D11463 7FC00297
@00000093 DB828293 00029103 00000013 00200113 00200E93 01300E13 01D11463
@0000009A 01C01A63 FF000513 00000593 00B52023 FF5FF06F FF000513 00100593
@000000A1 00B52023 FF5FF06F
