/* http://srecord.sourceforge.net/ */
@00000000 FF0100B7 F0008093 0F0F1137 F0F10113 0020C1B3 F00FFEB7 00FE8E93
@00000007 00200E13 4BD19063 0FF010B7 FF008093 F0F0F137 0F010113 0020C1B3
@0000000E FF010EB7 F00E8E93 00300E13 47D19E63 00FF00B7 0FF08093 0F0F1137
@00000015 F0F10113 0020C1B3 0FF01EB7 FF0E8E93 00400E13 45D19C63 F00FF0B7
@0000001C 00F08093 F0F0F137 0F010113 0020C1B3 00FF0EB7 0FFE8E93 00500E13
@00000023 43D19A63 FF0100B7 F0008093 0F0F1137 F0F10113 0020C0B3 F00FFEB7
@0000002A 00FE8E93 00600E13 41D09863 FF0100B7 F0008093 0F0F1137 F0F10113
@00000031 0020C133 F00FFEB7 00FE8E93 00700E13 3FD11663 FF0100B7 F0008093
@00000038 0010C0B3 00000E93 00800E13 3DD09A63 00000213 FF0100B7 F0008093
@0000003F 0F0F1137 F0F10113 0020C1B3 00018313 00120213 00200293 FE5210E3
@00000046 F00FFEB7 00FE8E93 00900E13 39D31E63 00000213 0FF010B7 FF008093
@0000004D F0F0F137 0F010113 0020C1B3 00000013 00018313 00120213 00200293
@00000054 FC521EE3 FF010EB7 F00E8E93 00A00E13 37D31063 00000213 00FF00B7
@0000005B 0FF08093 0F0F1137 F0F10113 0020C1B3 00000013 00000013 00018313
@00000062 00120213 00200293 FC521CE3 0FF01EB7 FF0E8E93 00B00E13 33D31063
@00000069 00000213 FF0100B7 F0008093 0F0F1137 F0F10113 0020C1B3 00120213
@00000070 00200293 FE5212E3 F00FFEB7 00FE8E93 00C00E13 2FD19663 00000213
@00000077 0FF010B7 FF008093 F0F0F137 0F010113 00000013 0020C1B3 00120213
@0000007E 00200293 FE5210E3 FF010EB7 F00E8E93 00D00E13 2BD19A63 00000213
@00000085 00FF00B7 0FF08093 0F0F1137 F0F10113 00000013 00000013 0020C1B3
@0000008C 00120213 00200293 FC521EE3 0FF01EB7 FF0E8E93 00E00E13 27D19C63
@00000093 00000213 FF0100B7 F0008093 00000013 0F0F1137 F0F10113 0020C1B3
@0000009A 00120213 00200293 FE5210E3 F00FFEB7 00FE8E93 00F00E13 25D19063
@000000A1 00000213 0FF010B7 FF008093 00000013 F0F0F137 0F010113 00000013
@000000A8 0020C1B3 00120213 00200293 FC521EE3 FF010EB7 F00E8E93 01000E13
@000000AF 21D19263 00000213 00FF00B7 0FF08093 00000013 00000013 0F0F1137
@000000B6 F0F10113 0020C1B3 00120213 00200293 FC521EE3 0FF01EB7 FF0E8E93
@000000BD 01100E13 1DD19463 00000213 0F0F1137 F0F10113 FF0100B7 F0008093
@000000C4 0020C1B3 00120213 00200293 FE5212E3 F00FFEB7 00FE8E93 01200E13
@000000CB 19D19A63 00000213 F0F0F137 0F010113 0FF010B7 FF008093 00000013
@000000D2 0020C1B3 00120213 00200293 FE5210E3 FF010EB7 F00E8E93 01300E13
@000000D9 15D19E63 00000213 0F0F1137 F0F10113 00FF00B7 0FF08093 00000013
@000000E0 00000013 0020C1B3 00120213 00200293 FC521EE3 0FF01EB7 FF0E8E93
@000000E7 01400E13 13D19063 00000213 0F0F1137 F0F10113 00000013 FF0100B7
@000000EE F0008093 0020C1B3 00120213 00200293 FE5210E3 F00FFEB7 00FE8E93
@000000F5 01500E13 0FD19463 00000213 F0F0F137 0F010113 00000013 0FF010B7
@000000FC FF008093 00000013 0020C1B3 00120213 00200293 FC521EE3 FF010EB7
@00000103 F00E8E93 01600E13 0BD19663 00000213 0F0F1137 F0F10113 00000013
@0000010A 00000013 00FF00B7 0FF08093 0020C1B3 00120213 00200293 FC521EE3
@00000111 0FF01EB7 FF0E8E93 01700E13 07D19863 FF0100B7 F0008093 00104133
@00000118 FF010EB7 F00E8E93 01800E13 05D11A63 00FF00B7 0FF08093 0000C133
@0000011F 00FF0EB7 0FFE8E93 01900E13 03D11C63 000040B3 00000E93 01A00E13
@00000126 03D09463 111110B7 11108093 22222137 22210113 0020C033 00000E93
@0000012D 01B00E13 01D01463 01C01A63 FF000513 00000593 00B52023 FF5FF06F
@00000134 FF000513 00100593 00B52023 FF5FF06F
