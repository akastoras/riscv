/* http://srecord.sourceforge.net/ */
@00000000 00FF10B7 F0008093 F0F0C193 FF00FEB7 00FE8E93 00200E13 1DD19663
@00000007 0FF010B7 FF008093 0F00C193 0FF01EB7 F00E8E93 00300E13 1BD19863
@0000000E 00FF10B7 8FF08093 70F0C193 00FF1EB7 FF0E8E93 00400E13 19D19A63
@00000015 F00FF0B7 00F08093 0F00C193 F00FFEB7 0FFE8E93 00500E13 17D19C63
@0000001C FF00F0B7 70008093 70F0C093 FF00FEB7 00FE8E93 00600E13 15D09E63
@00000023 00000213 0FF010B7 FF008093 0F00C193 00018313 00120213 00200293
@0000002A FE5214E3 0FF01EB7 F00E8E93 00700E13 13D31663 00000213 00FF10B7
@00000031 8FF08093 70F0C193 00000013 00018313 00120213 00200293 FE5212E3
@00000038 00FF1EB7 FF0E8E93 00800E13 0FD31C63 00000213 F00FF0B7 00F08093
@0000003F 0F00C193 00000013 00000013 00018313 00120213 00200293 FE5210E3
@00000046 F00FFEB7 0FFE8E93 00900E13 0DD31063 00000213 0FF010B7 FF008093
@0000004D 0F00C193 00120213 00200293 FE5216E3 0FF01EB7 F00E8E93 00A00E13
@00000054 09D19A63 00000213 00FF10B7 FFF08093 00000013 00F0C193 00120213
@0000005B 00200293 FE5214E3 00FF1EB7 FF0E8E93 00B00E13 07D19263 00000213
@00000062 F00FF0B7 00F08093 00000013 00000013 0F00C193 00120213 00200293
@00000069 FE5212E3 F00FFEB7 0FFE8E93 00C00E13 03D19863 0F004093 0F000E93
@00000070 00D00E13 03D09063 00FF00B7 0FF08093 70F0C013 00000E93 00E00E13
@00000077 01D01463 01C01A63 FF000513 00000593 00B52023 FF5FF06F FF000513
@0000007E 00100593 00B52023 FF5FF06F
