/* http://srecord.sourceforge.net/ */
@00000000 7FC00097 00008093 00008183 FFF00E93 00200E13 23D19C63 7FC00097
@00000007 FE808093 00108183 00000E93 00300E13 23D19063 7FC00097 FD008093
@0000000E 00208183 FF000E93 00400E13 21D19463 7FC00097 FB808093 00308183
@00000015 00F00E93 00500E13 1FD19863 7FC00097 FA308093 FFD08183 FFF00E93
@0000001C 00600E13 1DD19C63 7FC00097 F8B08093 FFE08183 00000E93 00700E13
@00000023 1DD19063 7FC00097 F7308093 FFF08183 FF000E93 00800E13 1BD19463
@0000002A 7FC00097 F5B08093 00008183 00F00E93 00900E13 19D19863 7FC00097
@00000031 F4008093 FE008093 02008283 FFF00E93 00A00E13 17D29A63 7FC00097
@00000038 F2408093 FFA08093 00708283 00000E93 00B00E13 15D29C63 00C00E13
@0000003F 00000213 7FC00097 F0108093 00108183 00018313 FF000E93 13D31C63
@00000046 00120213 00200293 FE5210E3 00D00E13 00000213 7FC00097 ED608093
@0000004D 00108183 00000013 00018313 00F00E93 11D31463 00120213 00200293
@00000054 FC521EE3 00E00E13 00000213 7FC00097 EA408093 00108183 00000013
@0000005B 00000013 00018313 00000E93 0DD31A63 00120213 00200293 FC521CE3
@00000062 00F00E13 00000213 7FC00097 E7108093 00108183 FF000E93 0BD19663
@00000069 00120213 00200293 FE5212E3 01000E13 00000213 7FC00097 E4A08093
@00000070 00000013 00108183 00F00E93 09D19063 00120213 00200293 FE5210E3
@00000077 01100E13 00000213 7FC00097 E1C08093 00000013 00000013 00108183
@0000007E 00000E93 05D19863 00120213 00200293 FC521EE3 7FC00297 DF428293
@00000085 00028103 00200113 00200E93 01200E13 03D11463 7FC00297 DD828293
@0000008C 00028103 00000013 00200113 00200E93 01300E13 01D11463 01C01A63
@00000093 FF000513 00000593 00B52023 FF5FF06F FF000513 00100593 00B52023
@0000009A FF5FF06F
