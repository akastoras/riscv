/* http://srecord.sourceforge.net/ */
@00000000 800000B7 0000D193 80000EB7 00200E13 29D19863 800000B7 0010D193
@00000007 40000EB7 00300E13 27D19E63 800000B7 0070D193 01000EB7 00400E13
@0000000E 27D19463 800000B7 00E0D193 00020EB7 00500E13 25D19A63 800000B7
@00000015 00108093 01F0D193 00100E93 00600E13 23D19E63 FFF00093 0000D193
@0000001C FFF00E93 00700E13 23D19463 FFF00093 0010D193 80000EB7 FFFE8E93
@00000023 00800E13 21D19863 FFF00093 0070D193 02000EB7 FFFE8E93 00900E13
@0000002A 1FD19C63 FFF00093 00E0D193 00040EB7 FFFE8E93 00A00E13 1FD19063
@00000031 FFF00093 01F0D193 00100E93 00B00E13 1DD19663 212120B7 12108093
@00000038 0000D193 21212EB7 121E8E93 00C00E13 1BD19863 212120B7 12108093
@0000003F 0010D193 10909EB7 090E8E93 00D00E13 19D19A63 212120B7 12108093
@00000046 0070D193 00424EB7 242E8E93 00E00E13 17D19C63 212120B7 12108093
@0000004D 00E0D193 00008EB7 484E8E93 00F00E13 15D19E63 212120B7 12108093
@00000054 01F0D193 00000E93 01000E13 15D19263 800000B7 0070D093 01000EB7
@0000005B 01100E13 13D09863 00000213 800000B7 0070D193 00018313 00120213
@00000062 00200293 FE5216E3 01000EB7 01200E13 11D31463 00000213 800000B7
@00000069 00E0D193 00000013 00018313 00120213 00200293 FE5214E3 00020EB7
@00000070 01300E13 0DD31E63 00000213 800000B7 00108093 01F0D193 00000013
@00000077 00000013 00018313 00120213 00200293 FE5210E3 00100E93 01400E13
@0000007E 0BD31463 00000213 800000B7 0070D193 00120213 00200293 FE5218E3
@00000085 01000EB7 01500E13 09D19263 00000213 800000B7 00000013 00E0D193
@0000008C 00120213 00200293 FE5216E3 00020EB7 01600E13 05D19E63 00000213
@00000093 800000B7 00108093 00000013 00000013 01F0D193 00120213 00200293
@0000009A FE5212E3 00100E93 01700E13 03D19663 00405093 00000E93 01800E13
@000000A1 01D09E63 02100093 00A0D013 00000E93 01900E13 01D01463 01C01A63
@000000A8 FF000513 00000593 00B52023 FF5FF06F FF000513 00100593 00B52023
@000000AF FF5FF06F
