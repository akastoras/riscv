/* http://srecord.sourceforge.net/ */
@00000000 7FC00097 00008093 00AA0137 0AA10113 0020A023 0000A183 00AA0EB7
@00000007 0AAE8E93 00200E13 47D19063 7FC00097 FD808093 AA00B137 A0010113
@0000000E 0020A223 0040A183 AA00BEB7 A00E8E93 00300E13 43D19C63 7FC00097
@00000015 FB008093 0AA01137 AA010113 0020A423 0080A183 0AA01EB7 AA0E8E93
@0000001C 00400E13 41D19863 7FC00097 F8808093 A00AA137 00A10113 0020A623
@00000023 00C0A183 A00AAEB7 00AE8E93 00500E13 3FD19463 7FC00097 F7C08093
@0000002A 00AA0137 0AA10113 FE20AA23 FF40A183 00AA0EB7 0AAE8E93 00600E13
@00000031 3DD19063 7FC00097 F5408093 AA00B137 A0010113 FE20AC23 FF80A183
@00000038 AA00BEB7 A00E8E93 00700E13 39D19C63 7FC00097 F2C08093 0AA01137
@0000003F AA010113 FE20AE23 FFC0A183 0AA01EB7 AA0E8E93 00800E13 37D19863
@00000046 7FC00097 F0408093 A00AA137 00A10113 0020A023 0000A183 A00AAEB7
@0000004D 00AE8E93 00900E13 35D19463 7FC00097 EE008093 12345137 67810113
@00000054 FE008213 02222023 0000A283 12345EB7 678E8E93 00A00E13 31D29E63
@0000005B 7FC00097 EB408093 58213137 09810113 FFD08093 0020A3A3 7FC00217
@00000062 EA020213 00022283 58213EB7 098E8E93 00B00E13 2FD29463 00C00E13
@00000069 00000213 AABBD0B7 CDD08093 7FC00117 E5010113 00112023 00012183
@00000070 AABBDEB7 CDDE8E93 2BD19E63 00120213 00200293 FC521AE3 00D00E13
@00000077 00000213 DAABC0B7 CCD08093 7FC00117 E1810113 00000013 00112223
@0000007E 00412183 DAABCEB7 CCDE8E93 29D19063 00120213 00200293 FC5218E3
@00000085 00E00E13 00000213 DDAAC0B7 BCC08093 7FC00117 DDC10113 00000013
@0000008C 00000013 00112423 00812183 DDAACEB7 BCCE8E93 25D19063 00120213
@00000093 00200293 FC5216E3 00F00E13 00000213 CDDAB0B7 BBC08093 00000013
@0000009A 7FC00117 D9810113 00112623 00C12183 CDDABEB7 BBCE8E93 21D19263
@000000A1 00120213 00200293 FC5218E3 01000E13 00000213 CCDDB0B7 ABB08093
@000000A8 00000013 7FC00117 D5C10113 00000013 00112823 01012183 CCDDBEB7
@000000AF ABBE8E93 1DD19263 00120213 00200293 FC5216E3 01100E13 00000213
@000000B6 BCCDE0B7 AAB08093 00000013 00000013 7FC00117 D1810113 00112A23
@000000BD 01412183 BCCDEEB7 AABE8E93 19D19263 00120213 00200293 FC5216E3
@000000C4 01200E13 00000213 7FC00117 CE810113 001120B7 23308093 00112023
@000000CB 00012183 00112EB7 233E8E93 15D19663 00120213 00200293 FC521AE3
@000000D2 01300E13 00000213 7FC00117 CB010113 300110B7 22308093 00000013
@000000D9 00112223 00412183 30011EB7 223E8E93 11D19863 00120213 00200293
@000000E0 FC5218E3 01400E13 00000213 7FC00117 C7410113 330010B7 12208093
@000000E7 00000013 00000013 00112423 00812183 33001EB7 122E8E93 0DD19863
@000000EE 00120213 00200293 FC5216E3 01500E13 00000213 7FC00117 C3410113
@000000F5 00000013 233000B7 11208093 00112623 00C12183 23300EB7 112E8E93
@000000FC 09D19A63 00120213 00200293 FC5218E3 01600E13 00000213 7FC00117
@00000103 BF810113 00000013 223300B7 01108093 00000013 00112823 01012183
@0000010A 22330EB7 011E8E93 05D19A63 00120213 00200293 FC5216E3 01700E13
@00000111 00000213 7FC00117 BB810113 00000013 00000013 122330B7 00108093
@00000118 00112A23 01412183 12233EB7 001E8E93 01D19A63 00120213 00200293
@0000011F FC5216E3 01C01A63 FF000513 00000593 00B52023 FF5FF06F FF000513
@00000126 00100593 00B52023 FF5FF06F
