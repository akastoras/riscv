/* http://srecord.sourceforge.net/ */
@00000000 7FC00097 00008093 0000D183 0FF00E93 00200E13 27D19663 7FC00097
@00000007 FE808093 0020D183 00010EB7 F00E8E93 00300E13 25D19863 7FC00097
@0000000E FCC08093 0040D183 00001EB7 FF0E8E93 00400E13 23D19A63 7FC00097
@00000015 FB008093 0060D183 0000FEB7 00FE8E93 00500E13 21D19C63 7FC00097
@0000001C F9A08093 FFA0D183 0FF00E93 00600E13 21D19063 7FC00097 F8208093
@00000023 FFC0D183 00010EB7 F00E8E93 00700E13 1FD19263 7FC00097 F6608093
@0000002A FFE0D183 00001EB7 FF0E8E93 00800E13 1DD19463 7FC00097 F4A08093
@00000031 0000D183 0000FEB7 00FE8E93 00900E13 1BD19663 7FC00097 F2808093
@00000038 FE008093 0200D283 0FF00E93 00A00E13 19D29863 7FC00097 F0C08093
@0000003F FFB08093 0070D283 00010EB7 F00E8E93 00B00E13 17D29863 00C00E13
@00000046 00000213 7FC00097 EE608093 0020D183 00018313 00001EB7 FF0E8E93
@0000004D 15D31663 00120213 00200293 FC521EE3 00D00E13 00000213 7FC00097
@00000054 EB808093 0020D183 00000013 00018313 0000FEB7 00FE8E93 11D31C63
@0000005B 00120213 00200293 FC521CE3 00E00E13 00000213 7FC00097 E8008093
@00000062 0020D183 00000013 00000013 00018313 00010EB7 F00E8E93 0FD31063
@00000069 00120213 00200293 FC521AE3 00F00E13 00000213 7FC00097 E4A08093
@00000070 0020D183 00001EB7 FF0E8E93 0BD19A63 00120213 00200293 FE5210E3
@00000077 01000E13 00000213 7FC00097 E2008093 00000013 0020D183 0000FEB7
@0000007E 00FE8E93 09D19263 00120213 00200293 FC521EE3 01100E13 00000213
@00000085 7FC00097 DEC08093 00000013 00000013 0020D183 00010EB7 F00E8E93
@0000008C 05D19863 00120213 00200293 FC521CE3 7FC00297 DC028293 0002D103
@00000093 00200113 00200E93 01200E13 03D11463 7FC00297 DA428293 0002D103
@0000009A 00000013 00200113 00200E93 01300E13 01D11463 01C01A63 FF000513
@000000A1 00000593 00B52023 FF5FF06F FF000513 00100593 00B52023 FF5FF06F
