/* http://srecord.sourceforge.net/ */
@00000000 00200E13 00000293 00000317 01030313 000302E7 0C00006F 00000317
@00000007 FFC30313 0A629A63 00400E13 00000213 00000317 01030313 000309E7
@0000000E 09C01E63 00120213 00200293 FE5214E3 00500E13 00000213 00000317
@00000015 01430313 00000013 000309E7 07C01A63 00120213 00200293 FE5212E3
@0000001C 00600E13 00000213 00000317 01830313 00000013 00000013 000309E7
@00000023 05C01463 00120213 00200293 FE5210E3 00100293 00000317 01C30313
@0000002A FFC30067 00128293 00128293 00128293 00128293 00128293 00128293
@00000031 00400E93 00700E13 01D29463 01C01A63 FF000513 00000593 00B52023
@00000038 FF5FF06F FF000513 00100593 00B52023 FF5FF06F
