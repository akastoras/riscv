/* http://srecord.sourceforge.net/ */
@00000000 00100093 00000113 002091B3 00100E93 00200E13 53D19E63 00100093
@00000007 00100113 002091B3 00200E93 00300E13 53D19263 00100093 00700113
@0000000E 002091B3 08000E93 00400E13 51D19663 00100093 00E00113 002091B3
@00000015 00004EB7 00500E13 4FD19A63 00100093 01F00113 002091B3 80000EB7
@0000001C 00600E13 4DD19E63 FFF00093 00000113 002091B3 FFF00E93 00700E13
@00000023 4DD19263 FFF00093 00100113 002091B3 FFE00E93 00800E13 4BD19663
@0000002A FFF00093 00700113 002091B3 F8000E93 00900E13 49D19A63 FFF00093
@00000031 00E00113 002091B3 FFFFCEB7 00A00E13 47D19E63 FFF00093 01F00113
@00000038 002091B3 80000EB7 00B00E13 47D19263 212120B7 12108093 00000113
@0000003F 002091B3 21212EB7 121E8E93 00C00E13 45D19263 212120B7 12108093
@00000046 00100113 002091B3 42424EB7 242E8E93 00D00E13 43D19263 212120B7
@0000004D 12108093 00700113 002091B3 90909EB7 080E8E93 00E00E13 41D19263
@00000054 212120B7 12108093 00E00113 002091B3 48484EB7 00F00E13 3FD19463
@0000005B 212120B7 12108093 01F00113 002091B3 80000EB7 01000E13 3DD19663
@00000062 212120B7 12108093 FC000113 002091B3 21212EB7 121E8E93 01100E13
@00000069 3BD19663 212120B7 12108093 FC100113 002091B3 42424EB7 242E8E93
@00000070 01200E13 39D19663 212120B7 12108093 FC700113 002091B3 90909EB7
@00000077 080E8E93 01300E13 37D19663 212120B7 12108093 FCE00113 002091B3
@0000007E 48484EB7 01400E13 35D19863 00100093 00700113 002090B3 08000E93
@00000085 01600E13 33D09C63 00100093 00E00113 00209133 00004EB7 01700E13
@0000008C 33D11063 00300093 001090B3 01800E93 01800E13 31D09663 00000213
@00000093 00100093 00700113 002091B3 00018313 00120213 00200293 FE5214E3
@0000009A 08000E93 01900E13 2FD31063 00000213 00100093 00E00113 002091B3
@000000A1 00000013 00018313 00120213 00200293 FE5212E3 00004EB7 01A00E13
@000000A8 2BD31863 00000213 00100093 01F00113 002091B3 00000013 00000013
@000000AF 00018313 00120213 00200293 FE5210E3 80000EB7 01B00E13 27D31E63
@000000B6 00000213 00100093 00700113 002091B3 00120213 00200293 FE5216E3
@000000BD 08000E93 01C00E13 25D19A63 00000213 00100093 00E00113 00000013
@000000C4 002091B3 00120213 00200293 FE5214E3 00004EB7 01D00E13 23D19463
@000000CB 00000213 00100093 01F00113 00000013 00000013 002091B3 00120213
@000000D2 00200293 FE5212E3 80000EB7 01E00E13 1FD19C63 00000213 00100093
@000000D9 00000013 00700113 002091B3 00120213 00200293 FE5214E3 08000E93
@000000E0 01F00E13 1DD19663 00000213 00100093 00000013 00E00113 00000013
@000000E7 002091B3 00120213 00200293 FE5212E3 00004EB7 02000E13 19D19E63
@000000EE 00000213 00100093 00000013 00000013 01F00113 002091B3 00120213
@000000F5 00200293 FE5212E3 80000EB7 02100E13 17D19663 00000213 00700113
@000000FC 00100093 002091B3 00120213 00200293 FE5216E3 08000E93 02200E13
@00000103 15D19263 00000213 00E00113 00100093 00000013 002091B3 00120213
@0000010A 00200293 FE5214E3 00004EB7 02300E13 11D19C63 00000213 01F00113
@00000111 00100093 00000013 00000013 002091B3 00120213 00200293 FE5212E3
@00000118 80000EB7 02400E13 0FD19463 00000213 00700113 00000013 00100093
@0000011F 002091B3 00120213 00200293 FE5214E3 08000E93 02500E13 0BD19E63
@00000126 00000213 00E00113 00000013 00100093 00000013 002091B3 00120213
@0000012D 00200293 FE5212E3 00004EB7 02600E13 09D19663 00000213 01F00113
@00000134 00000013 00000013 00100093 002091B3 00120213 00200293 FE5212E3
@0000013B 80000EB7 02700E13 05D19E63 00F00093 00101133 00000E93 02800E13
@00000142 05D11463 02000093 00009133 02000E93 02900E13 03D11A63 000010B3
@00000149 00000E93 02A00E13 03D09263 40000093 00001137 80010113 00209033
@00000150 00000E93 02B00E13 01D01463 01C01A63 FF000513 00000593 00B52023
@00000157 FF5FF06F FF000513 00100593 00B52023 FF5FF06F
