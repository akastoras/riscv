/* http://srecord.sourceforge.net/ */
@00000000 FF0100B7 F0008093 F0F0F193 FF010EB7 F00E8E93 00200E13 1BD19463
@00000007 0FF010B7 FF008093 0F00F193 0F000E93 00300E13 19D19863 00FF00B7
@0000000E 0FF08093 70F0F193 00F00E93 00400E13 17D19C63 F00FF0B7 00F08093
@00000015 0F00F193 00000E93 00500E13 17D19063 FF0100B7 F0008093 0F00F093
@0000001C 00000E93 00600E13 15D09463 00000213 0FF010B7 FF008093 70F0F193
@00000023 00018313 00120213 00200293 FE5214E3 70000E93 00700E13 11D31E63
@0000002A 00000213 00FF00B7 0FF08093 0F00F193 00000013 00018313 00120213
@00000031 00200293 FE5212E3 0F000E93 00800E13 0FD31663 00000213 F00FF0B7
@00000038 00F08093 F0F0F193 00000013 00000013 00018313 00120213 00200293
@0000003F FE5210E3 F00FFEB7 00FE8E93 00900E13 0BD31A63 00000213 0FF010B7
@00000046 FF008093 70F0F193 00120213 00200293 FE5216E3 70000E93 00A00E13
@0000004D 09D19663 00000213 00FF00B7 0FF08093 00000013 0F00F193 00120213
@00000054 00200293 FE5214E3 0F000E93 00B00E13 07D19063 00000213 F00FF0B7
@0000005B 00F08093 00000013 00000013 70F0F193 00120213 00200293 FE5212E3
@00000062 00F00E93 00C00E13 03D19863 0F007093 00000E93 00D00E13 03D09063
@00000069 00FF00B7 0FF08093 70F0F013 00000E93 00E00E13 01D01463 01C01A63
@00000070 FF000513 00000593 00B52023 FF5FF06F FF000513 00100593 00B52023
@00000077 FF5FF06F
