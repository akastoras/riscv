/* http://srecord.sourceforge.net/ */
@00000000 7FC00097 00008093 0000A183 00FF0EB7 0FFE8E93 00200E13 27D19A63
@00000007 7FC00097 FE408093 0040A183 FF010EB7 F00E8E93 00300E13 25D19C63
@0000000E 7FC00097 FC808093 0080A183 0FF01EB7 FF0E8E93 00400E13 23D19E63
@00000015 7FC00097 FAC08093 00C0A183 F00FFEB7 00FE8E93 00500E13 23D19063
@0000001C 7FC00097 F9C08093 FF40A183 00FF0EB7 0FFE8E93 00600E13 21D19263
@00000023 7FC00097 F8008093 FF80A183 FF010EB7 F00E8E93 00700E13 1FD19463
@0000002A 7FC00097 F6408093 FFC0A183 0FF01EB7 FF0E8E93 00800E13 1DD19663
@00000031 7FC00097 F4808093 0000A183 F00FFEB7 00FE8E93 00900E13 1BD19863
@00000038 7FC00097 F2008093 FE008093 0200A283 00FF0EB7 0FFE8E93 00A00E13
@0000003F 19D29863 7FC00097 F0008093 FFD08093 0070A283 FF010EB7 F00E8E93
@00000046 00B00E13 17D29863 00C00E13 00000213 7FC00097 EDC08093 0040A183
@0000004D 00018313 0FF01EB7 FF0E8E93 15D31663 00120213 00200293 FC521EE3
@00000054 00D00E13 00000213 7FC00097 EB008093 0040A183 00000013 00018313
@0000005B F00FFEB7 00FE8E93 11D31C63 00120213 00200293 FC521CE3 00E00E13
@00000062 00000213 7FC00097 E7408093 0040A183 00000013 00000013 00018313
@00000069 FF010EB7 F00E8E93 0FD31063 00120213 00200293 FC521AE3 00F00E13
@00000070 00000213 7FC00097 E4008093 0040A183 0FF01EB7 FF0E8E93 0BD19A63
@00000077 00120213 00200293 FE5210E3 01000E13 00000213 7FC00097 E1808093
@0000007E 00000013 0040A183 F00FFEB7 00FE8E93 09D19263 00120213 00200293
@00000085 FC521EE3 01100E13 00000213 7FC00097 DE008093 00000013 00000013
@0000008C 0040A183 FF010EB7 F00E8E93 05D19863 00120213 00200293 FC521CE3
@00000093 7FC00297 DB428293 0002A103 00200113 00200E93 01200E13 03D11463
@0000009A 7FC00297 D9828293 0002A103 00000013 00200113 00200E93 01300E13
@000000A1 01D11463 01C01A63 FF000513 00000593 00B52023 FF5FF06F FF000513
@000000A8 00100593 00B52023 FF5FF06F
