/* http://srecord.sourceforge.net/ */
@00000000 800000B7 00000113 4020D1B3 80000EB7 00200E13 59D19463 800000B7
@00000007 00100113 4020D1B3 C0000EB7 00300E13 57D19863 800000B7 00700113
@0000000E 4020D1B3 FF000EB7 00400E13 55D19C63 800000B7 00E00113 4020D1B3
@00000015 FFFE0EB7 00500E13 55D19063 800000B7 00108093 01F00113 4020D1B3
@0000001C FFF00E93 00600E13 53D19263 800000B7 FFF08093 00000113 4020D1B3
@00000023 80000EB7 FFFE8E93 00700E13 51D19263 800000B7 FFF08093 00100113
@0000002A 4020D1B3 40000EB7 FFFE8E93 00800E13 4FD19263 800000B7 FFF08093
@00000031 00700113 4020D1B3 01000EB7 FFFE8E93 00900E13 4DD19263 800000B7
@00000038 FFF08093 00E00113 4020D1B3 00020EB7 FFFE8E93 00A00E13 4BD19263
@0000003F 800000B7 FFF08093 01F00113 4020D1B3 00000E93 00B00E13 49D19463
@00000046 818180B7 18108093 00000113 4020D1B3 81818EB7 181E8E93 00C00E13
@0000004D 47D19463 818180B7 18108093 00100113 4020D1B3 C0C0CEB7 0C0E8E93
@00000054 00D00E13 45D19463 818180B7 18108093 00700113 4020D1B3 FF030EB7
@0000005B 303E8E93 00E00E13 43D19463 818180B7 18108093 00E00113 4020D1B3
@00000062 FFFE0EB7 606E8E93 00F00E13 41D19463 818180B7 18108093 01F00113
@00000069 4020D1B3 FFF00E93 01000E13 3FD19663 818180B7 18108093 FC000113
@00000070 4020D1B3 81818EB7 181E8E93 01100E13 3DD19663 818180B7 18108093
@00000077 FC100113 4020D1B3 C0C0CEB7 0C0E8E93 01200E13 3BD19663 818180B7
@0000007E 18108093 FC700113 4020D1B3 FF030EB7 303E8E93 01300E13 39D19663
@00000085 818180B7 18108093 FCE00113 4020D1B3 FFFE0EB7 606E8E93 01400E13
@0000008C 37D19663 818180B7 18108093 FFF00113 4020D1B3 FFF00E93 01500E13
@00000093 35D19863 800000B7 00700113 4020D0B3 FF000EB7 01600E13 33D09C63
@0000009A 800000B7 00E00113 4020D133 FFFE0EB7 01700E13 33D11063 00700093
@000000A1 4010D0B3 00000E93 01800E13 31D09663 00000213 800000B7 00700113
@000000A8 4020D1B3 00018313 00120213 00200293 FE5214E3 FF000EB7 01900E13
@000000AF 2FD31063 00000213 800000B7 00E00113 4020D1B3 00000013 00018313
@000000B6 00120213 00200293 FE5212E3 FFFE0EB7 01A00E13 2BD31863 00000213
@000000BD 800000B7 01F00113 4020D1B3 00000013 00000013 00018313 00120213
@000000C4 00200293 FE5210E3 FFF00E93 01B00E13 27D31E63 00000213 800000B7
@000000CB 00700113 4020D1B3 00120213 00200293 FE5216E3 FF000EB7 01C00E13
@000000D2 25D19A63 00000213 800000B7 00E00113 00000013 4020D1B3 00120213
@000000D9 00200293 FE5214E3 FFFE0EB7 01D00E13 23D19463 00000213 800000B7
@000000E0 01F00113 00000013 00000013 4020D1B3 00120213 00200293 FE5212E3
@000000E7 FFF00E93 01E00E13 1FD19C63 00000213 800000B7 00000013 00700113
@000000EE 4020D1B3 00120213 00200293 FE5214E3 FF000EB7 01F00E13 1DD19663
@000000F5 00000213 800000B7 00000013 00E00113 00000013 4020D1B3 00120213
@000000FC 00200293 FE5212E3 FFFE0EB7 02000E13 19D19E63 00000213 800000B7
@00000103 00000013 00000013 01F00113 4020D1B3 00120213 00200293 FE5212E3
@0000010A FFF00E93 02100E13 17D19663 00000213 00700113 800000B7 4020D1B3
@00000111 00120213 00200293 FE5216E3 FF000EB7 02200E13 15D19263 00000213
@00000118 00E00113 800000B7 00000013 4020D1B3 00120213 00200293 FE5214E3
@0000011F FFFE0EB7 02300E13 11D19C63 00000213 01F00113 800000B7 00000013
@00000126 00000013 4020D1B3 00120213 00200293 FE5212E3 FFF00E93 02400E13
@0000012D 0FD19463 00000213 00700113 00000013 800000B7 4020D1B3 00120213
@00000134 00200293 FE5214E3 FF000EB7 02500E13 0BD19E63 00000213 00E00113
@0000013B 00000013 800000B7 00000013 4020D1B3 00120213 00200293 FE5212E3
@00000142 FFFE0EB7 02600E13 09D19663 00000213 01F00113 00000013 00000013
@00000149 800000B7 4020D1B3 00120213 00200293 FE5212E3 FFF00E93 02700E13
@00000150 05D19E63 00F00093 40105133 00000E93 02800E13 05D11463 02000093
@00000157 4000D133 02000E93 02900E13 03D11A63 400050B3 00000E93 02A00E13
@0000015E 03D09263 40000093 00001137 80010113 4020D033 00000E93 02B00E13
@00000165 01D01463 01C01A63 FF000513 00000593 00B52023 FF5FF06F FF000513
@0000016C 00100593 00B52023 FF5FF06F
