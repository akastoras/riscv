/* http://srecord.sourceforge.net/ */
@00000000 00200E13 00000093 00000113 0020D663 31C01863 01C01663 FE20DEE3
@00000007 31C01263 00300E13 00100093 00100113 0020D663 2FC01863 01C01663
@0000000E FE20DEE3 2FC01263 00400E13 FFF00093 FFF00113 0020D663 2DC01863
@00000015 01C01663 FE20DEE3 2DC01263 00500E13 00100093 00000113 0020D663
@0000001C 2BC01863 01C01663 FE20DEE3 2BC01263 00600E13 00100093 FFF00113
@00000023 0020D663 29C01863 01C01663 FE20DEE3 29C01263 00700E13 FFF00093
@0000002A FFE00113 0020D663 27C01863 01C01663 FE20DEE3 27C01263 00800E13
@00000031 00000093 00100113 0020D463 01C01463 25C01663 FE20DEE3 00900E13
@00000038 FFF00093 00100113 0020D463 01C01463 23C01863 FE20DEE3 00A00E13
@0000003F FFE00093 FFF00113 0020D463 01C01463 21C01A63 FE20DEE3 00B00E13
@00000046 FFE00093 00100113 0020D463 01C01463 1FC01C63 FE20DEE3 00C00E13
@0000004D 00000213 FFF00093 00000113 1E20D063 00120213 00200293 FE5216E3
@00000054 00D00E13 00000213 FFF00093 00000113 00000013 1A20DE63 00120213
@0000005B 00200293 FE5214E3 00E00E13 00000213 FFF00093 00000113 00000013
@00000062 00000013 1820DA63 00120213 00200293 FE5212E3 00F00E13 00000213
@00000069 FFF00093 00000013 00000113 1620D863 00120213 00200293 FE5214E3
@00000070 01000E13 00000213 FFF00093 00000013 00000113 00000013 1420D463
@00000077 00120213 00200293 FE5212E3 01100E13 00000213 FFF00093 00000013
@0000007E 00000013 00000113 1220D063 00120213 00200293 FE5212E3 01200E13
@00000085 00000213 FFF00093 00000113 1020D063 00120213 00200293 FE5216E3
@0000008C 01300E13 00000213 FFF00093 00000113 00000013 0C20DE63 00120213
@00000093 00200293 FE5214E3 01400E13 00000213 FFF00093 00000113 00000013
@0000009A 00000013 0A20DA63 00120213 00200293 FE5212E3 01500E13 00000213
@000000A1 FFF00093 00000013 00000113 0820D863 00120213 00200293 FE5214E3
@000000A8 01600E13 00000213 FFF00093 00000013 00000113 00000013 0620D463
@000000AF 00120213 00200293 FE5212E3 01700E13 00000213 FFF00093 00000013
@000000B6 00000013 00000113 0420D063 00120213 00200293 FE5212E3 00100093
@000000BD 0000DA63 00108093 00108093 00108093 00108093 00108093 00108093
@000000C4 00300E93 01800E13 01D09463 01C01A63 FF000513 00000593 00B52023
@000000CB FF5FF06F FF000513 00100593 00B52023 FF5FF06F
