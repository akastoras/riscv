/* http://srecord.sourceforge.net/ */
@00000000 FF0100B7 F0008093 F0F0E193 F0F00E93 00200E13 1DD19463 0FF010B7
@00000007 FF008093 0F00E193 0FF01EB7 FF0E8E93 00300E13 1BD19663 00FF00B7
@0000000E 0FF08093 70F0E193 00FF0EB7 7FFE8E93 00400E13 19D19863 F00FF0B7
@00000015 00F08093 0F00E193 F00FFEB7 0FFE8E93 00500E13 17D19A63 FF0100B7
@0000001C F0008093 0F00E093 FF010EB7 FF0E8E93 00600E13 15D09C63 00000213
@00000023 0FF010B7 FF008093 0F00E193 00018313 00120213 00200293 FE5214E3
@0000002A 0FF01EB7 FF0E8E93 00700E13 13D31463 00000213 00FF00B7 0FF08093
@00000031 70F0E193 00000013 00018313 00120213 00200293 FE5212E3 00FF0EB7
@00000038 7FFE8E93 00800E13 0FD31A63 00000213 F00FF0B7 00F08093 0F00E193
@0000003F 00000013 00000013 00018313 00120213 00200293 FE5210E3 F00FFEB7
@00000046 0FFE8E93 00900E13 0BD31E63 00000213 0FF010B7 FF008093 0F00E193
@0000004D 00120213 00200293 FE5216E3 0FF01EB7 FF0E8E93 00A00E13 09D19863
@00000054 00000213 00FF00B7 0FF08093 00000013 F0F0E193 00120213 00200293
@0000005B FE5214E3 FFF00E93 00B00E13 07D19263 00000213 F00FF0B7 00F08093
@00000062 00000013 00000013 0F00E193 00120213 00200293 FE5212E3 F00FFEB7
@00000069 0FFE8E93 00C00E13 03D19863 0F006093 0F000E93 00D00E13 03D09063
@00000070 00FF00B7 0FF08093 70F0E013 00000E93 00E00E13 01D01463 01C01A63
@00000077 FF000513 00000593 00B52023 FF5FF06F FF000513 00100593 00B52023
@0000007E FF5FF06F
