/* http://srecord.sourceforge.net/ */
@00000000 00200E13 00000093 00100113 00209663 2BC01A63 01C01663 FE209EE3
@00000007 2BC01463 00300E13 00100093 00000113 00209663 29C01A63 01C01663
@0000000E FE209EE3 29C01463 00400E13 FFF00093 00100113 00209663 27C01A63
@00000015 01C01663 FE209EE3 27C01463 00500E13 00100093 FFF00113 00209663
@0000001C 25C01A63 01C01663 FE209EE3 25C01463 00600E13 00000093 00000113
@00000023 00209463 01C01463 23C01863 FE209EE3 00700E13 00100093 00100113
@0000002A 00209463 01C01463 21C01A63 FE209EE3 00800E13 FFF00093 FFF00113
@00000031 00209463 01C01463 1FC01C63 FE209EE3 00900E13 00000213 00000093
@00000038 00000113 1E209063 00120213 00200293 FE5216E3 00A00E13 00000213
@0000003F 00000093 00000113 00000013 1A209E63 00120213 00200293 FE5214E3
@00000046 00B00E13 00000213 00000093 00000113 00000013 00000013 18209A63
@0000004D 00120213 00200293 FE5212E3 00C00E13 00000213 00000093 00000013
@00000054 00000113 16209863 00120213 00200293 FE5214E3 00D00E13 00000213
@0000005B 00000093 00000013 00000113 00000013 14209463 00120213 00200293
@00000062 FE5212E3 00E00E13 00000213 00000093 00000013 00000013 00000113
@00000069 12209063 00120213 00200293 FE5212E3 00F00E13 00000213 00000093
@00000070 00000113 10209063 00120213 00200293 FE5216E3 01000E13 00000213
@00000077 00000093 00000113 00000013 0C209E63 00120213 00200293 FE5214E3
@0000007E 01100E13 00000213 00000093 00000113 00000013 00000013 0A209A63
@00000085 00120213 00200293 FE5212E3 01200E13 00000213 00000093 00000013
@0000008C 00000113 08209863 00120213 00200293 FE5214E3 01300E13 00000213
@00000093 00000093 00000013 00000113 00000013 06209463 00120213 00200293
@0000009A FE5212E3 01400E13 00000213 00000093 00000013 00000013 00000113
@000000A1 04209063 00120213 00200293 FE5212E3 00100093 00009A63 00108093
@000000A8 00108093 00108093 00108093 00108093 00108093 00300E93 01500E13
@000000AF 01D09463 01C01A63 FF000513 00000593 00B52023 FF5FF06F FF000513
@000000B6 00100593 00B52023 FF5FF06F
