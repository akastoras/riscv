/* http://srecord.sourceforge.net/ */
@00000000 00000093 4000D193 00000E93 00200E13 2BD19463 800000B7 4010D193
@00000007 C0000EB7 00300E13 29D19A63 800000B7 4070D193 FF000EB7 00400E13
@0000000E 29D19063 800000B7 40E0D193 FFFE0EB7 00500E13 27D19663 800000B7
@00000015 00108093 41F0D193 FFF00E93 00600E13 25D19A63 800000B7 FFF08093
@0000001C 4000D193 80000EB7 FFFE8E93 00700E13 23D19C63 800000B7 FFF08093
@00000023 4010D193 40000EB7 FFFE8E93 00800E13 21D19E63 800000B7 FFF08093
@0000002A 4070D193 01000EB7 FFFE8E93 00900E13 21D19063 800000B7 FFF08093
@00000031 40E0D193 00020EB7 FFFE8E93 00A00E13 1FD19263 800000B7 FFF08093
@00000038 41F0D193 00000E93 00B00E13 1DD19663 818180B7 18108093 4000D193
@0000003F 81818EB7 181E8E93 00C00E13 1BD19863 818180B7 18108093 4010D193
@00000046 C0C0CEB7 0C0E8E93 00D00E13 19D19A63 818180B7 18108093 4070D193
@0000004D FF030EB7 303E8E93 00E00E13 17D19C63 818180B7 18108093 40E0D193
@00000054 FFFE0EB7 606E8E93 00F00E13 15D19E63 818180B7 18108093 41F0D193
@0000005B FFF00E93 01000E13 15D19263 800000B7 4070D093 FF000EB7 01100E13
@00000062 13D09863 00000213 800000B7 4070D193 00018313 00120213 00200293
@00000069 FE5216E3 FF000EB7 01200E13 11D31463 00000213 800000B7 40E0D193
@00000070 00000013 00018313 00120213 00200293 FE5214E3 FFFE0EB7 01300E13
@00000077 0DD31E63 00000213 800000B7 00108093 41F0D193 00000013 00000013
@0000007E 00018313 00120213 00200293 FE5210E3 FFF00E93 01400E13 0BD31463
@00000085 00000213 800000B7 4070D193 00120213 00200293 FE5218E3 FF000EB7
@0000008C 01500E13 09D19263 00000213 800000B7 00000013 40E0D193 00120213
@00000093 00200293 FE5216E3 FFFE0EB7 01600E13 05D19E63 00000213 800000B7
@0000009A 00108093 00000013 00000013 41F0D193 00120213 00200293 FE5212E3
@000000A1 FFF00E93 01700E13 03D19663 40405093 00000E93 01800E13 01D09E63
@000000A8 02100093 40A0D013 00000E93 01900E13 01D01463 01C01A63 FF000513
@000000AF 00000593 00B52023 FF5FF06F FF000513 00100593 00B52023 FF5FF06F
