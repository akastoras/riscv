/* http://srecord.sourceforge.net/ */
@00000000 00000093 0000A193 00000E93 00200E13 27D19263 00100093 0010A193
@00000007 00000E93 00300E13 25D19863 00300093 0070A193 00100E93 00400E13
@0000000E 23D19E63 00700093 0030A193 00000E93 00500E13 23D19463 00000093
@00000015 8000A193 00000E93 00600E13 21D19A63 800000B7 0000A193 00100E93
@0000001C 00700E13 21D19063 800000B7 8000A193 00100E93 00800E13 1FD19663
@00000023 00000093 7FF0A193 00100E93 00900E13 1DD19C63 800000B7 FFF08093
@0000002A 0000A193 00000E93 00A00E13 1DD19063 800000B7 FFF08093 7FF0A193
@00000031 00000E93 00B00E13 1BD19463 800000B7 7FF0A193 00100E93 00C00E13
@00000038 19D19A63 800000B7 FFF08093 8000A193 00000E93 00D00E13 17D19E63
@0000003F 00000093 FFF0A193 00000E93 00E00E13 17D19463 FFF00093 0010A193
@00000046 00100E93 00F00E13 15D19A63 FFF00093 FFF0A193 00000E93 01000E13
@0000004D 15D19063 00B00093 00D0A093 00100E93 01100E13 13D09663 00000213
@00000054 00F00093 00A0A193 00018313 00120213 00200293 FE5216E3 00000E93
@0000005B 01200E13 11D31263 00000213 00A00093 0100A193 00000013 00018313
@00000062 00120213 00200293 FE5214E3 00100E93 01300E13 0DD31C63 00000213
@00000069 01000093 0090A193 00000013 00000013 00018313 00120213 00200293
@00000070 FE5212E3 00000E93 01400E13 0BD31463 00000213 00B00093 00F0A193
@00000077 00120213 00200293 FE5218E3 00100E93 01500E13 09D19263 00000213
@0000007E 01100093 00000013 0080A193 00120213 00200293 FE5216E3 00000E93
@00000085 01600E13 05D19E63 00000213 00C00093 00000013 00000013 00E0A193
@0000008C 00120213 00200293 FE5214E3 00100E93 01700E13 03D19863 FFF02093
@00000093 00000E93 01800E13 03D09063 00FF00B7 0FF08093 FFF0A013 00000E93
@0000009A 01900E13 01D01463 01C01A63 FF000513 00000593 00B52023 FF5FF06F
@000000A1 FF000513 00100593 00B52023 FF5FF06F
