/* http://srecord.sourceforge.net/ */
@00000000 800000B7 00000113 0020D1B3 80000EB7 00200E13 57D19863 800000B7
@00000007 00100113 0020D1B3 40000EB7 00300E13 55D19C63 800000B7 00700113
@0000000E 0020D1B3 01000EB7 00400E13 55D19063 800000B7 00E00113 0020D1B3
@00000015 00020EB7 00500E13 53D19463 800000B7 00108093 01F00113 0020D1B3
@0000001C 00100E93 00600E13 51D19663 FFF00093 00000113 0020D1B3 FFF00E93
@00000023 00700E13 4FD19A63 FFF00093 00100113 0020D1B3 80000EB7 FFFE8E93
@0000002A 00800E13 4DD19C63 FFF00093 00700113 0020D1B3 02000EB7 FFFE8E93
@00000031 00900E13 4BD19E63 FFF00093 00E00113 0020D1B3 00040EB7 FFFE8E93
@00000038 00A00E13 4BD19063 FFF00093 01F00113 0020D1B3 00100E93 00B00E13
@0000003F 49D19463 212120B7 12108093 00000113 0020D1B3 21212EB7 121E8E93
@00000046 00C00E13 47D19463 212120B7 12108093 00100113 0020D1B3 10909EB7
@0000004D 090E8E93 00D00E13 45D19463 212120B7 12108093 00700113 0020D1B3
@00000054 00424EB7 242E8E93 00E00E13 43D19463 212120B7 12108093 00E00113
@0000005B 0020D1B3 00008EB7 484E8E93 00F00E13 41D19463 212120B7 12108093
@00000062 01F00113 0020D1B3 00000E93 01000E13 3FD19663 212120B7 12108093
@00000069 FC000113 0020D1B3 21212EB7 121E8E93 01100E13 3DD19663 212120B7
@00000070 12108093 FC100113 0020D1B3 10909EB7 090E8E93 01200E13 3BD19663
@00000077 212120B7 12108093 FC700113 0020D1B3 00424EB7 242E8E93 01300E13
@0000007E 39D19663 212120B7 12108093 FCE00113 0020D1B3 00008EB7 484E8E93
@00000085 01400E13 37D19663 212120B7 12108093 FFF00113 0020D1B3 00000E93
@0000008C 01500E13 35D19863 800000B7 00700113 0020D0B3 01000EB7 01600E13
@00000093 33D09C63 800000B7 00E00113 0020D133 00020EB7 01700E13 33D11063
@0000009A 00700093 0010D0B3 00000E93 01800E13 31D09663 00000213 800000B7
@000000A1 00700113 0020D1B3 00018313 00120213 00200293 FE5214E3 01000EB7
@000000A8 01900E13 2FD31063 00000213 800000B7 00E00113 0020D1B3 00000013
@000000AF 00018313 00120213 00200293 FE5212E3 00020EB7 01A00E13 2BD31863
@000000B6 00000213 800000B7 01F00113 0020D1B3 00000013 00000013 00018313
@000000BD 00120213 00200293 FE5210E3 00100E93 01B00E13 27D31E63 00000213
@000000C4 800000B7 00700113 0020D1B3 00120213 00200293 FE5216E3 01000EB7
@000000CB 01C00E13 25D19A63 00000213 800000B7 00E00113 00000013 0020D1B3
@000000D2 00120213 00200293 FE5214E3 00020EB7 01D00E13 23D19463 00000213
@000000D9 800000B7 01F00113 00000013 00000013 0020D1B3 00120213 00200293
@000000E0 FE5212E3 00100E93 01E00E13 1FD19C63 00000213 800000B7 00000013
@000000E7 00700113 0020D1B3 00120213 00200293 FE5214E3 01000EB7 01F00E13
@000000EE 1DD19663 00000213 800000B7 00000013 00E00113 00000013 0020D1B3
@000000F5 00120213 00200293 FE5212E3 00020EB7 02000E13 19D19E63 00000213
@000000FC 800000B7 00000013 00000013 01F00113 0020D1B3 00120213 00200293
@00000103 FE5212E3 00100E93 02100E13 17D19663 00000213 00700113 800000B7
@0000010A 0020D1B3 00120213 00200293 FE5216E3 01000EB7 02200E13 15D19263
@00000111 00000213 00E00113 800000B7 00000013 0020D1B3 00120213 00200293
@00000118 FE5214E3 00020EB7 02300E13 11D19C63 00000213 01F00113 800000B7
@0000011F 00000013 00000013 0020D1B3 00120213 00200293 FE5212E3 00100E93
@00000126 02400E13 0FD19463 00000213 00700113 00000013 800000B7 0020D1B3
@0000012D 00120213 00200293 FE5214E3 01000EB7 02500E13 0BD19E63 00000213
@00000134 00E00113 00000013 800000B7 00000013 0020D1B3 00120213 00200293
@0000013B FE5212E3 00020EB7 02600E13 09D19663 00000213 01F00113 00000013
@00000142 00000013 800000B7 0020D1B3 00120213 00200293 FE5212E3 00100E93
@00000149 02700E13 05D19E63 00F00093 00105133 00000E93 02800E13 05D11463
@00000150 02000093 0000D133 02000E93 02900E13 03D11A63 000050B3 00000E93
@00000157 02A00E13 03D09263 40000093 00001137 80010113 0020D033 00000E93
@0000015E 02B00E13 01D01463 01C01A63 FF000513 00000593 00B52023 FF5FF06F
@00000165 FF000513 00100593 00B52023 FF5FF06F
