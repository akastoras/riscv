/* http://srecord.sourceforge.net/ */
@00000000 00000093 00000113 402081B3 00000E93 00200E13 4BD19663 00100093
@00000007 00100113 402081B3 00000E93 00300E13 49D19A63 00300093 00700113
@0000000E 402081B3 FFC00E93 00400E13 47D19E63 00000093 FFFF8137 402081B3
@00000015 00008EB7 00500E13 47D19263 800000B7 00000113 402081B3 80000EB7
@0000001C 00600E13 45D19663 800000B7 FFFF8137 402081B3 80008EB7 00700E13
@00000023 43D19A63 00000093 00008137 FFF10113 402081B3 FFFF8EB7 001E8E93
@0000002A 00800E13 41D19A63 800000B7 FFF08093 00000113 402081B3 80000EB7
@00000031 FFFE8E93 00900E13 3FD19A63 800000B7 FFF08093 00008137 FFF10113
@00000038 402081B3 7FFF8EB7 00A00E13 3DD19A63 800000B7 00008137 FFF10113
@0000003F 402081B3 7FFF8EB7 001E8E93 00B00E13 3BD19A63 800000B7 FFF08093
@00000046 FFFF8137 402081B3 80008EB7 FFFE8E93 00C00E13 39D19A63 00000093
@0000004D FFF00113 402081B3 00100E93 00D00E13 37D19E63 FFF00093 00100113
@00000054 402081B3 FFE00E93 00E00E13 37D19263 FFF00093 FFF00113 402081B3
@0000005B 00000E93 00F00E13 35D19663 00D00093 00B00113 402080B3 00200E93
@00000062 01000E13 33D09A63 00E00093 00B00113 40208133 00300E93 01100E13
@00000069 31D11E63 00D00093 401080B3 00000E93 01200E13 31D09463 00000213
@00000070 00D00093 00B00113 402081B3 00018313 00120213 00200293 FE5214E3
@00000077 00200E93 01300E13 2DD31E63 00000213 00E00093 00B00113 402081B3
@0000007E 00000013 00018313 00120213 00200293 FE5212E3 00300E93 01400E13
@00000085 2BD31663 00000213 00F00093 00B00113 402081B3 00000013 00000013
@0000008C 00018313 00120213 00200293 FE5210E3 00400E93 01500E13 27D31C63
@00000093 00000213 00D00093 00B00113 402081B3 00120213 00200293 FE5216E3
@0000009A 00200E93 01600E13 25D19863 00000213 00E00093 00B00113 00000013
@000000A1 402081B3 00120213 00200293 FE5214E3 00300E93 01700E13 23D19263
@000000A8 00000213 00F00093 00B00113 00000013 00000013 402081B3 00120213
@000000AF 00200293 FE5212E3 00400E93 01800E13 1FD19A63 00000213 00D00093
@000000B6 00000013 00B00113 402081B3 00120213 00200293 FE5214E3 00200E93
@000000BD 01900E13 1DD19463 00000213 00E00093 00000013 00B00113 00000013
@000000C4 402081B3 00120213 00200293 FE5212E3 00300E93 01A00E13 19D19C63
@000000CB 00000213 00F00093 00000013 00000013 00B00113 402081B3 00120213
@000000D2 00200293 FE5212E3 00400E93 01B00E13 17D19463 00000213 00B00113
@000000D9 00D00093 402081B3 00120213 00200293 FE5216E3 00200E93 01C00E13
@000000E0 15D19063 00000213 00B00113 00E00093 00000013 402081B3 00120213
@000000E7 00200293 FE5214E3 00300E93 01D00E13 11D19A63 00000213 00B00113
@000000EE 00F00093 00000013 00000013 402081B3 00120213 00200293 FE5212E3
@000000F5 00400E93 01E00E13 0FD19263 00000213 00B00113 00000013 00D00093
@000000FC 402081B3 00120213 00200293 FE5214E3 00200E93 01F00E13 0BD19C63
@00000103 00000213 00B00113 00000013 00E00093 00000013 402081B3 00120213
@0000010A 00200293 FE5212E3 00300E93 02000E13 09D19463 00000213 00B00113
@00000111 00000013 00000013 00F00093 402081B3 00120213 00200293 FE5212E3
@00000118 00400E93 02100E13 05D19C63 FF100093 40100133 00F00E93 02200E13
@0000011F 05D11263 02000093 40008133 02000E93 02300E13 03D11863 400000B3
@00000126 00000E93 02400E13 03D09063 01000093 01E00113 40208033 00000E93
@0000012D 02500E13 01D01463 01C01A63 FF000513 00000593 00B52023 FF5FF06F
@00000134 FF000513 00100593 00B52023 FF5FF06F
