/* http://srecord.sourceforge.net/ */
@00000000 00200E13 00000093 00100113 0020E663 2FC01263 01C01663 FE20EEE3
@00000007 2DC01C63 00300E13 FFE00093 FFF00113 0020E663 2DC01263 01C01663
@0000000E FE20EEE3 2BC01C63 00400E13 00000093 FFF00113 0020E663 2BC01263
@00000015 01C01663 FE20EEE3 29C01C63 00500E13 00100093 00000113 0020E463
@0000001C 01C01463 29C01063 FE20EEE3 00600E13 FFF00093 FFE00113 0020E463
@00000023 01C01463 27C01263 FE20EEE3 00700E13 FFF00093 00000113 0020E463
@0000002A 01C01463 25C01463 FE20EEE3 00800E13 800000B7 80000137 FFF10113
@00000031 0020E463 01C01463 23C01463 FE20EEE3 00900E13 00000213 F00000B7
@00000038 F0000137 FFF10113 2020E663 00120213 00200293 FE5214E3 00A00E13
@0000003F 00000213 F00000B7 F0000137 FFF10113 00000013 1E20E263 00120213
@00000046 00200293 FE5212E3 00B00E13 00000213 F00000B7 F0000137 FFF10113
@0000004D 00000013 00000013 1A20EC63 00120213 00200293 FE5210E3 00C00E13
@00000054 00000213 F00000B7 00000013 F0000137 FFF10113 1820E863 00120213
@0000005B 00200293 FE5212E3 00D00E13 00000213 F00000B7 00000013 F0000137
@00000062 FFF10113 00000013 1620E263 00120213 00200293 FE5210E3 00E00E13
@00000069 00000213 F00000B7 00000013 00000013 F0000137 FFF10113 1220EC63
@00000070 00120213 00200293 FE5210E3 00F00E13 00000213 F00000B7 F0000137
@00000077 FFF10113 1020EA63 00120213 00200293 FE5214E3 01000E13 00000213
@0000007E F00000B7 F0000137 FFF10113 00000013 0E20E663 00120213 00200293
@00000085 FE5212E3 01100E13 00000213 F00000B7 F0000137 FFF10113 00000013
@0000008C 00000013 0C20E063 00120213 00200293 FE5210E3 01200E13 00000213
@00000093 F00000B7 00000013 F0000137 FFF10113 0820EC63 00120213 00200293
@0000009A FE5212E3 01300E13 00000213 F00000B7 00000013 F0000137 FFF10113
@000000A1 00000013 0620E663 00120213 00200293 FE5210E3 01400E13 00000213
@000000A8 F00000B7 00000013 00000013 F0000137 FFF10113 0420E063 00120213
@000000AF 00200293 FE5210E3 00100093 00106A63 00108093 00108093 00108093
@000000B6 00108093 00108093 00108093 00300E93 01500E13 01D09463 01C01A63
@000000BD FF000513 00000593 00B52023 FF5FF06F FF000513 00100593 00B52023
@000000C4 FF5FF06F
