/* http://srecord.sourceforge.net/ */
@00000000 7FC00097 00008093 FAA00113 00208023 00008183 FAA00E93 00200E13
@00000007 3DD19C63 7FC00097 FE008093 00000113 002080A3 00108183 00000E93
@0000000E 00300E13 3BD19C63 7FC00097 FC008093 FFFFF137 FA010113 00208123
@00000015 00209183 FFFFFEB7 FA0E8E93 00400E13 39D19863 7FC00097 F9808093
@0000001C 00A00113 002081A3 00308183 00A00E93 00500E13 37D19863 7FC00097
@00000023 F7F08093 FAA00113 FE208EA3 FFD08183 FAA00E93 00600E13 35D19863
@0000002A 7FC00097 F5F08093 00000113 FE208F23 FFE08183 00000E93 00700E13
@00000031 33D19863 7FC00097 F3F08093 FA000113 FE208FA3 FFF08183 FA000E93
@00000038 00800E13 31D19863 7FC00097 F1F08093 00A00113 00208023 00008183
@0000003F 00A00E93 00900E13 2FD19863 7FC00097 F0008093 12345137 67810113
@00000046 FE008213 02220023 00008283 07800E93 00A00E13 2DD29463 7FC00097
@0000004D ED808093 00003137 09810113 FFA08093 002083A3 7FC00217 EC120213
@00000054 00020283 F9800E93 00B00E13 29D29C63 00C00E13 00000213 FDD00093
@0000005B 7FC00117 E9410113 00110023 00010183 FDD00E93 27D19A63 00120213
@00000062 00200293 FC521EE3 00D00E13 00000213 FCD00093 7FC00117 E6410113
@00000069 00000013 001100A3 00110183 FCD00E93 25D19063 00120213 00200293
@00000070 FC521CE3 00E00E13 00000213 FCC00093 7FC00117 E3010113 00000013
@00000077 00000013 00110123 00210183 FCC00E93 21D19463 00120213 00200293
@0000007E FC521AE3 00F00E13 00000213 FBC00093 00000013 7FC00117 DF410113
@00000085 001101A3 00310183 FBC00E93 1DD19A63 00120213 00200293 FC521CE3
@0000008C 01000E13 00000213 FBB00093 00000013 7FC00117 DC010113 00000013
@00000093 00110223 00410183 FBB00E93 19D19E63 00120213 00200293 FC521AE3
@0000009A 01100E13 00000213 FAB00093 00000013 00000013 7FC00117 D8410113
@000000A1 001102A3 00510183 FAB00E93 17D19263 00120213 00200293 FC521AE3
@000000A8 01200E13 00000213 7FC00117 D5810113 03300093 00110023 00010183
@000000AF 03300E93 13D19A63 00120213 00200293 FC521EE3 01300E13 00000213
@000000B6 7FC00117 D2810113 02300093 00000013 001100A3 00110183 02300E93
@000000BD 11D19063 00120213 00200293 FC521CE3 01400E13 00000213 7FC00117
@000000C4 CF410113 02200093 00000013 00000013 00110123 00210183 02200E93
@000000CB 0DD19463 00120213 00200293 FC521AE3 01500E13 00000213 7FC00117
@000000D2 CBC10113 00000013 01200093 001101A3 00310183 01200E93 09D19A63
@000000D9 00120213 00200293 FC521CE3 01600E13 00000213 7FC00117 C8810113
@000000E0 00000013 01100093 00000013 00110223 00410183 01100E93 05D19E63
@000000E7 00120213 00200293 FC521AE3 01700E13 00000213 7FC00117 C5010113
@000000EE 00000013 00000013 00100093 001102A3 00510183 00100E93 03D19263
@000000F5 00120213 00200293 FC521AE3 0EF00513 7FC00597 C1C58593 00A581A3
@000000FC 01C01A63 FF000513 00000593 00B52023 FF5FF06F FF000513 00100593
@00000103 00B52023 FF5FF06F
