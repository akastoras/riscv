/* http://srecord.sourceforge.net/ */
@00000000 00100093 00009193 00100E93 00200E13 27D19A63 00100093 00109193
@00000007 00200E93 00300E13 27D19063 00100093 00709193 08000E93 00400E13
@0000000E 25D19663 00100093 00E09193 00004EB7 00500E13 23D19C63 00100093
@00000015 01F09193 80000EB7 00600E13 23D19263 FFF00093 00009193 FFF00E93
@0000001C 00700E13 21D19863 FFF00093 00109193 FFE00E93 00800E13 1FD19E63
@00000023 FFF00093 00709193 F8000E93 00900E13 1FD19463 FFF00093 00E09193
@0000002A FFFFCEB7 00A00E13 1DD19A63 FFF00093 01F09193 80000EB7 00B00E13
@00000031 1DD19063 212120B7 12108093 00009193 21212EB7 121E8E93 00C00E13
@00000038 1BD19263 212120B7 12108093 00109193 42424EB7 242E8E93 00D00E13
@0000003F 19D19463 212120B7 12108093 00709193 90909EB7 080E8E93 00E00E13
@00000046 17D19663 212120B7 12108093 00E09193 48484EB7 00F00E13 15D19A63
@0000004D 212120B7 12108093 01F09193 80000EB7 01000E13 13D19E63 00100093
@00000054 00709093 08000E93 01100E13 13D09463 00000213 00100093 00709193
@0000005B 00018313 00120213 00200293 FE5216E3 08000E93 01200E13 11D31063
@00000062 00000213 00100093 00E09193 00000013 00018313 00120213 00200293
@00000069 FE5214E3 00004EB7 01300E13 0DD31A63 00000213 00100093 01F09193
@00000070 00000013 00000013 00018313 00120213 00200293 FE5212E3 80000EB7
@00000077 01400E13 0BD31263 00000213 00100093 00709193 00120213 00200293
@0000007E FE5218E3 08000E93 01500E13 09D19063 00000213 00100093 00000013
@00000085 00E09193 00120213 00200293 FE5216E3 00004EB7 01600E13 05D19C63
@0000008C 00000213 00100093 00000013 00000013 01F09193 00120213 00200293
@00000093 FE5214E3 80000EB7 01700E13 03D19663 01F01093 00000E93 01800E13
@0000009A 01D09E63 02100093 01409013 00000E93 01900E13 01D01463 01C01A63
@000000A1 FF000513 00000593 00B52023 FF5FF06F FF000513 00100593 00B52023
@000000A8 FF5FF06F
