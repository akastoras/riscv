/* http://srecord.sourceforge.net/ */
@00000000 7FC00097 00008093 0AA00113 00209023 00009183 0AA00E93 00200E13
@00000007 45D19E63 7FC00097 FE008093 FFFFB137 A0010113 00209123 00209183
@0000000E FFFFBEB7 A00E8E93 00300E13 43D19A63 7FC00097 FB808093 BEEF1137
@00000015 AA010113 00209223 0040A183 BEEF1EB7 AA0E8E93 00400E13 41D19663
@0000001C 7FC00097 F9008093 FFFFA137 00A10113 00209323 00609183 FFFFAEB7
@00000023 00AE8E93 00500E13 3FD19263 7FC00097 F7608093 0AA00113 FE209D23
@0000002A FFA09183 0AA00E93 00600E13 3DD19263 7FC00097 F5608093 FFFFB137
@00000031 A0010113 FE209E23 FFC09183 FFFFBEB7 A00E8E93 00700E13 39D19E63
@00000038 7FC00097 F2E08093 00001137 AA010113 FE209F23 FFE09183 00001EB7
@0000003F AA0E8E93 00800E13 37D19A63 7FC00097 F0608093 FFFFA137 00A10113
@00000046 00209023 00009183 FFFFAEB7 00AE8E93 00900E13 35D19663 7FC00097
@0000004D EE008093 12345137 67810113 FE008213 02221023 00009283 00005EB7
@00000054 678E8E93 00A00E13 33D29063 7FC00097 EB408093 00003137 09810113
@0000005B FFB08093 002093A3 7FC00217 E9E20213 00021283 00003EB7 098E8E93
@00000062 00B00E13 2FD29663 00C00E13 00000213 FFFFD0B7 CDD08093 7FC00117
@00000069 E6010113 00111023 00011183 FFFFDEB7 CDDE8E93 2DD19063 00120213
@00000070 00200293 FC521AE3 00D00E13 00000213 FFFFC0B7 CCD08093 7FC00117
@00000077 E2810113 00000013 00111123 00211183 FFFFCEB7 CCDE8E93 29D19263
@0000007E 00120213 00200293 FC5218E3 00E00E13 00000213 FFFFC0B7 BCC08093
@00000085 7FC00117 DEC10113 00000013 00000013 00111223 00411183 FFFFCEB7
@0000008C BCCE8E93 25D19263 00120213 00200293 FC5216E3 00F00E13 00000213
@00000093 FFFFB0B7 BBC08093 00000013 7FC00117 DA810113 00111323 00611183
@0000009A FFFFBEB7 BBCE8E93 21D19463 00120213 00200293 FC5218E3 01000E13
@000000A1 00000213 FFFFB0B7 ABB08093 00000013 7FC00117 D6C10113 00000013
@000000A8 00111423 00811183 FFFFBEB7 ABBE8E93 1DD19463 00120213 00200293
@000000AF FC5216E3 01100E13 00000213 FFFFE0B7 AAB08093 00000013 00000013
@000000B6 7FC00117 D2810113 00111523 00A11183 FFFFEEB7 AABE8E93 19D19463
@000000BD 00120213 00200293 FC5216E3 01200E13 00000213 7FC00117 CF810113
@000000C4 000020B7 23308093 00111023 00011183 00002EB7 233E8E93 15D19863
@000000CB 00120213 00200293 FC521AE3 01300E13 00000213 7FC00117 CC010113
@000000D2 000010B7 22308093 00000013 00111123 00211183 00001EB7 223E8E93
@000000D9 11D19A63 00120213 00200293 FC5218E3 01400E13 00000213 7FC00117
@000000E0 C8410113 000010B7 12208093 00000013 00000013 00111223 00411183
@000000E7 00001EB7 122E8E93 0DD19A63 00120213 00200293 FC5216E3 01500E13
@000000EE 00000213 7FC00117 C4410113 00000013 11200093 00111323 00611183
@000000F5 11200E93 0BD19063 00120213 00200293 FC521CE3 01600E13 00000213
@000000FC 7FC00117 C1010113 00000013 01100093 00000013 00111423 00811183
@00000103 01100E93 07D19463 00120213 00200293 FC521AE3 01700E13 00000213
@0000010A 7FC00117 BD810113 00000013 00000013 000030B7 00108093 00111523
@00000111 00A11183 00003EB7 001E8E93 03D19463 00120213 00200293 FC5216E3
@00000118 0000C537 EEF50513 7FC00597 B9858593 00A59323 01C01A63 FF000513
@0000011F 00000593 00B52023 FF5FF06F FF000513 00100593 00B52023 FF5FF06F
