/* http://srecord.sourceforge.net/ */
@00000000 FF0100B7 F0008093 0F0F1137 F0F10113 0020E1B3 FF100EB7 F0FE8E93
@00000007 00200E13 4BD19263 0FF010B7 FF008093 F0F0F137 0F010113 0020E1B3
@0000000E FFF10EB7 FF0E8E93 00300E13 49D19063 00FF00B7 0FF08093 0F0F1137
@00000015 F0F10113 0020E1B3 0FFF1EB7 FFFE8E93 00400E13 45D19E63 F00FF0B7
@0000001C 00F08093 F0F0F137 0F010113 0020E1B3 F0FFFEB7 0FFE8E93 00500E13
@00000023 43D19C63 FF0100B7 F0008093 0F0F1137 F0F10113 0020E0B3 FF100EB7
@0000002A F0FE8E93 00600E13 41D09A63 FF0100B7 F0008093 0F0F1137 F0F10113
@00000031 0020E133 FF100EB7 F0FE8E93 00700E13 3FD11863 FF0100B7 F0008093
@00000038 0010E0B3 FF010EB7 F00E8E93 00800E13 3DD09A63 00000213 FF0100B7
@0000003F F0008093 0F0F1137 F0F10113 0020E1B3 00018313 00120213 00200293
@00000046 FE5210E3 FF100EB7 F0FE8E93 00900E13 39D31E63 00000213 0FF010B7
@0000004D FF008093 F0F0F137 0F010113 0020E1B3 00000013 00018313 00120213
@00000054 00200293 FC521EE3 FFF10EB7 FF0E8E93 00A00E13 37D31063 00000213
@0000005B 00FF00B7 0FF08093 0F0F1137 F0F10113 0020E1B3 00000013 00000013
@00000062 00018313 00120213 00200293 FC521CE3 0FFF1EB7 FFFE8E93 00B00E13
@00000069 33D31063 00000213 FF0100B7 F0008093 0F0F1137 F0F10113 0020E1B3
@00000070 00120213 00200293 FE5212E3 FF100EB7 F0FE8E93 00C00E13 2FD19663
@00000077 00000213 0FF010B7 FF008093 F0F0F137 0F010113 00000013 0020E1B3
@0000007E 00120213 00200293 FE5210E3 FFF10EB7 FF0E8E93 00D00E13 2BD19A63
@00000085 00000213 00FF00B7 0FF08093 0F0F1137 F0F10113 00000013 00000013
@0000008C 0020E1B3 00120213 00200293 FC521EE3 0FFF1EB7 FFFE8E93 00E00E13
@00000093 27D19C63 00000213 FF0100B7 F0008093 00000013 0F0F1137 F0F10113
@0000009A 0020E1B3 00120213 00200293 FE5210E3 FF100EB7 F0FE8E93 00F00E13
@000000A1 25D19063 00000213 0FF010B7 FF008093 00000013 F0F0F137 0F010113
@000000A8 00000013 0020E1B3 00120213 00200293 FC521EE3 FFF10EB7 FF0E8E93
@000000AF 01000E13 21D19263 00000213 00FF00B7 0FF08093 00000013 00000013
@000000B6 0F0F1137 F0F10113 0020E1B3 00120213 00200293 FC521EE3 0FFF1EB7
@000000BD FFFE8E93 01100E13 1DD19463 00000213 0F0F1137 F0F10113 FF0100B7
@000000C4 F0008093 0020E1B3 00120213 00200293 FE5212E3 FF100EB7 F0FE8E93
@000000CB 01200E13 19D19A63 00000213 F0F0F137 0F010113 0FF010B7 FF008093
@000000D2 00000013 0020E1B3 00120213 00200293 FE5210E3 FFF10EB7 FF0E8E93
@000000D9 01300E13 15D19E63 00000213 0F0F1137 F0F10113 00FF00B7 0FF08093
@000000E0 00000013 00000013 0020E1B3 00120213 00200293 FC521EE3 0FFF1EB7
@000000E7 FFFE8E93 01400E13 13D19063 00000213 0F0F1137 F0F10113 00000013
@000000EE FF0100B7 F0008093 0020E1B3 00120213 00200293 FE5210E3 FF100EB7
@000000F5 F0FE8E93 01500E13 0FD19463 00000213 F0F0F137 0F010113 00000013
@000000FC 0FF010B7 FF008093 00000013 0020E1B3 00120213 00200293 FC521EE3
@00000103 FFF10EB7 FF0E8E93 01600E13 0BD19663 00000213 0F0F1137 F0F10113
@0000010A 00000013 00000013 00FF00B7 0FF08093 0020E1B3 00120213 00200293
@00000111 FC521EE3 0FFF1EB7 FFFE8E93 01700E13 07D19863 FF0100B7 F0008093
@00000118 00106133 FF010EB7 F00E8E93 01800E13 05D11A63 00FF00B7 0FF08093
@0000011F 0000E133 00FF0EB7 0FFE8E93 01900E13 03D11C63 000060B3 00000E93
@00000126 01A00E13 03D09463 111110B7 11108093 22222137 22210113 0020E033
@0000012D 00000E93 01B00E13 01D01463 01C01A63 FF000513 00000593 00B52023
@00000134 FF5FF06F FF000513 00100593 00B52023 FF5FF06F
