/* http://srecord.sourceforge.net/ */
@00000000 00002517 71C50513 004005EF 40B50533 00002EB7 710E8E93 00200E13
@00000007 03D51463 FFFFE517 8FC50513 004005EF 40B50533 FFFFEEB7 8F0E8E93
@0000000E 00300E13 01D51463 01C01A63 FF000513 00000593 00B52023 FF5FF06F
@00000015 FF000513 00100593 00B52023 FF5FF06F 00000000
