/* http://srecord.sourceforge.net/ */
@00000000 00000093 00008193 00000E93 00200E13 27D19C63 00100093 00108193
@00000007 00200E93 00300E13 27D19263 00300093 00708193 00A00E93 00400E13
@0000000E 25D19863 00000093 80008193 80000E93 00500E13 23D19E63 800000B7
@00000015 00008193 80000EB7 00600E13 23D19463 800000B7 80008193 80000EB7
@0000001C 800E8E93 00700E13 21D19863 00000093 7FF08193 7FF00E93 00800E13
@00000023 1FD19E63 800000B7 FFF08093 00008193 80000EB7 FFFE8E93 00900E13
@0000002A 1FD19063 800000B7 FFF08093 7FF08193 80000EB7 7FEE8E93 00A00E13
@00000031 1DD19263 800000B7 7FF08193 80000EB7 7FFE8E93 00B00E13 1BD19663
@00000038 800000B7 FFF08093 80008193 7FFFFEB7 7FFE8E93 00C00E13 19D19863
@0000003F 00000093 FFF08193 FFF00E93 00D00E13 17D19E63 FFF00093 00108193
@00000046 00000E93 00E00E13 17D19463 FFF00093 FFF08193 FFE00E93 00F00E13
@0000004D 15D19A63 800000B7 FFF08093 00108193 80000EB7 01000E13 13D19E63
@00000054 00D00093 00B08093 01800E93 01100E13 13D09463 00000213 00D00093
@0000005B 00B08193 00018313 00120213 00200293 FE5216E3 01800E93 01200E13
@00000062 11D31063 00000213 00D00093 00A08193 00000013 00018313 00120213
@00000069 00200293 FE5214E3 01700E93 01300E13 0DD31A63 00000213 00D00093
@00000070 00908193 00000013 00000013 00018313 00120213 00200293 FE5212E3
@00000077 01600E93 01400E13 0BD31263 00000213 00D00093 00B08193 00120213
@0000007E 00200293 FE5218E3 01800E93 01500E13 09D19063 00000213 00D00093
@00000085 00000013 00A08193 00120213 00200293 FE5216E3 01700E93 01600E13
@0000008C 05D19C63 00000213 00D00093 00000013 00000013 00908193 00120213
@00000093 00200293 FE5214E3 01600E93 01700E13 03D19663 02000093 02000E93
@0000009A 01800E13 01D09E63 02100093 03208013 00000E93 01900E13 01D01463
@000000A1 01C01A63 FF000513 00000593 00B52023 FF5FF06F FF000513 00100593
@000000A8 00B52023 FF5FF06F
